/*module alu(
    input [31:0] A, B,
    input [1:0] ALUOp,
    output [31:0] ALUResult
);

always @ (*)
begin
    casex (ALUOp)
        00:
        01:
        10:
 
        default: 
    endcase
end*/

aa
